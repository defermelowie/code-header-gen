----------------------------------------------------------
-- Test project
----------------------------------------------------------
-- A project to test sgen
--
-- File: test.vhd (vhdl)
-- By: Lowie Deferme (UHasselt/KULeuven - FIIW)
-- On: 02 February 2022